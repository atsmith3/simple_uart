
`ifndef __DATATYPES_SV__
`define __DATATYPES_SV__

typedef enum bit [8:0] {
  B_4800=96,
  B_9600=48,
  B_19200=24,
  B_38400=12,
  B_57600=8,
  B_115200=4,
} baud_t;

`endif
